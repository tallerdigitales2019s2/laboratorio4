module TecTacToe();

endmodule