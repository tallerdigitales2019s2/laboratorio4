//module Game(clk, btn_right_i, btn_down_i, btn_confirm_i,board_status_o,current_scrren_o,current_player_o);
//endmodule