module TecTacToe();
endmodule